`ifndef SUM
`define SUM

module sum(
    input [15:0] a,
    input [15:0] b,
    output [15:0] result
);

    assign result = a + b;
endmodule
`endif
